`include "CONFIG_MACROS_SYS.v"
module system_top (
    input   wire    REF_CLK,
    input   wire    UART_CLK,
    input   wire    RST,
    input   wire    RX_IN,
    output  wire    TX_OUT
);
////////////////////////////////////////////////////////////////////////////////
/////////////////////// internal wires of RegFile /////////////////////////////
//////////////////////////////////////////////////////////////////////////////
wire    WrEn_top,
        SYNC_RST_REF_CLK,
        RdEn_top,
        RdData_VLD_top;

wire    [`ADDR-1:0]     Address_top;

wire    [`WIDTH-1:0]    WrData_top,
                        RdData_top,
                        REG0_OP_A,
                        REG1_OP_B,
                        REG2_UART_convig,
                        REG3_div ;
///////////////////////////////////////////////////////////////////////////////
///////////////////////////// internal wires of ALU //////////////////////////
/////////////////////////////////////////////////////////////////////////////
wire    EN_top,
        ALU_CLK,
        OUT_VALID_top;

wire    [3:0]   ALU_FUN_top;

wire    [`WIDTH_OUT_ALU-1:0]    ALU_OUT_top;
////////////////////////////////////////////////////////////////////////////////
//////////////////////////// internal wires of UART ///////////////////////////
//////////////////////////////////////////////////////////////////////////////
wire  [`WIDTH-1:0]  TX_IN_DATA_top,
                    RX_out_DATA_top;

wire  TX_IN_valid_top,
      CLK_TX_top,
      SYNC_RST_UART_CLK,
      TX_busy,
      RX_out_valid_top;

wire  I_clk_en_top;

wire  Gate_EN;

wire  [`WIDTH-1:0]  sync_RX_OUT_DATA;
wire  sync_RX_OUT_V;

wire  [`WIDTH-1:0]  CTRL_out_DATA;
wire  CTRL_out_V;

wire  SYNC_TX_busy;
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////// SYS_CTRL ////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
SYS_CTRL U0_CTRL_TOP(
    //CTRL_RX
    .UART_RX_DATA(sync_RX_OUT_DATA),
    .UART_RX_VLD(sync_RX_OUT_V),
    .CLK(REF_CLK),
    .RST(SYNC_RST_REF_CLK),
    .ALU_EN(EN_top),
    .ALU_FUN(ALU_FUN_top),
    .CLKG_EN(Gate_EN),
    .RF_Address(Address_top),
    .RF_WrEn(WrEn_top),
    .RF_RdEn(RdEn_top),
    .RF_WrData(WrData_top),
    //CTRL_TX
    .ALU_OUT(ALU_OUT_top),
    .ALU_OUT_VLD(OUT_VALID_top),
    .RF_RdData(RdData_top),
    .RF_RdData_VLD(RdData_VLD_top),
    .UART_TX_Busy(TX_busy),
    .UART_TX_DATA(CTRL_out_DATA),
    .UART_TX_VLD(CTRL_out_V),
    .CLKDIV_EN(I_clk_en_top)
);
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////// RegFile ////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
RegFile UO_RegFile(
.CLK(REF_CLK),
.RST(SYNC_RST_REF_CLK),
.WrEn(WrEn_top),
.RdEn(RdEn_top),
.Address(Address_top),
.WrData(WrData_top),
.RdData(RdData_top),
.RdData_VLD(RdData_VLD_top),
.REG0(REG0_OP_A),
.REG1(REG1_OP_B),
.REG2(REG2_UART_convig),
.REG3(REG3_div)
);
////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////// ALU //////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
ALU U0_ALU
(
  .A(REG0_OP_A), 
  .B(REG1_OP_B),
  .EN(EN_top),
  .ALU_FUN(ALU_FUN_top),
  .CLK(ALU_CLK),
  .RST(SYNC_RST_REF_CLK),  
  .ALU_OUT(ALU_OUT_top),
  .OUT_VALID(OUT_VALID_top)  
);
////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////// UART /////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
UART_TOP U0_UART(
    .TX_IN_DATA(TX_IN_DATA_top),
    .RX_IN_DATA(RX_IN),
    .TX_IN_valid(TX_IN_valid_top),
    .CLK_RX(UART_CLK),
    .CLK_TX(CLK_TX_top),
    .parity_enable(REG2_UART_convig[0]),
    .RST(SYNC_RST_UART_CLK),
    .parity_type(REG2_UART_convig[1]),
    .prescale(REG2_UART_convig[6:2]),
    .TX_out_valid(TX_busy),
    .RX_out_valid(RX_out_valid_top),
    .TX_out_DATA(TX_OUT),
    .RX_out_DATA(RX_out_DATA_top)
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// clock divider ///////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
clock_divider U0_clock_divider(
  .I_div_ratio(REG3_div[4:0]),     ////////////////////////////////////////
  .I_ref_clk(UART_CLK),
  .I_clk_en(I_clk_en_top),
  .I_rst_n(SYNC_RST_UART_CLK),
  .o_div_clk(CLK_TX_top) 
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// clock Gating ///////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
CLK_GATE U0_CLK_GATE (
.CLK_EN(Gate_EN),
.CLK(REF_CLK),
.GATED_CLK(ALU_CLK)
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// Data Sync of RX /////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
data_synchronizer U0_Data_Sync_of_RX (
    .unsync_bus(RX_out_DATA_top),
    .bus_enable(RX_out_valid_top),
    .clk(REF_CLK),
    .rst(SYNC_RST_REF_CLK),
    .sync_bus(sync_RX_OUT_DATA),
    .enable_pulse(sync_RX_OUT_V)  
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// Data Sync of TX /////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
data_synchronizer U0_Data_Sync_of_TX (
    .unsync_bus(CTRL_out_DATA),
    .bus_enable(CTRL_out_V),
    .clk(CLK_TX_top),
    .rst(SYNC_RST_UART_CLK),
    .sync_bus(TX_IN_DATA_top),
    .enable_pulse(TX_IN_valid_top)  
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// SYNC RST UART CLK ///////////////////////////////
//////////////////////////////////////////////////////////////////////////////
RST_synchronizer U0_SYNC_RST_UART_CLK (
    .RST(RST),
    .clk(UART_CLK),
    .SYNC_RST(SYNC_RST_UART_CLK)
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// SYNC RST REF CLK ///////////////////////////////
//////////////////////////////////////////////////////////////////////////////
RST_synchronizer U0_SYNC_RST_REF_CLK (
    .RST(RST),
    .clk(REF_CLK),
    .SYNC_RST(SYNC_RST_REF_CLK)
);
////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////// SYNC Bit //////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
bit_synchronizer U0_bit_synchronizer (
    .ASYNC(TX_busy),
    .RST(SYNC_RST_REF_CLK),
    .clk(REF_CLK),
    .SYNC(SYNC_TX_busy)
);
endmodule
