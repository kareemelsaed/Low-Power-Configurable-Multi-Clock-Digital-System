`include "CONFIG_MACROS_SYS.v"
module system_top (
    input   wire    REF_CLK,
    input   wire    UART_CLK,
    input   wire    RST,
    input   wire    RX_IN,
/////////////////////////////////// DFT /////////////////////////////////
    input   wire  [`NUM_OF_CHAINS-1:0]  SI,
    input   wire                        SE,
    input   wire                        test_mode,
    input   wire                        scan_clk,
    input   wire                        scan_rst,
    output  wire  [`NUM_OF_CHAINS-1:0]  SO,
/////////////////////////////////////////////////////////////////////////
    output  wire    TX_OUT
);
////////////////////////////////////////////////////////////////////////////////
/////////////////////// internal wires of RegFile /////////////////////////////
//////////////////////////////////////////////////////////////////////////////
wire    WrEn_top,
        SYNC_RST_REF_CLK,
        RdEn_top,
        RdData_VLD_top;

wire    [`ADDR-1:0]     Address_top;

wire    [`WIDTH-1:0]    WrData_top,
                        RdData_top,
                        REG0_OP_A,
                        REG1_OP_B,
                        REG2_UART_convig,
                        REG3_div ;
///////////////////////////////////////////////////////////////////////////////
///////////////////////////// internal wires of ALU //////////////////////////
/////////////////////////////////////////////////////////////////////////////
wire    EN_top,
        ALU_CLK,
        OUT_VALID_top;

wire    [3:0]   ALU_FUN_top;

wire    [`WIDTH_OUT_ALU-1:0]    ALU_OUT_top;
////////////////////////////////////////////////////////////////////////////////
//////////////////////////// internal wires of UART ///////////////////////////
//////////////////////////////////////////////////////////////////////////////
wire  [`WIDTH-1:0]  TX_IN_DATA_top,
                    RX_out_DATA_top;

wire  TX_IN_valid_top,
      CLK_TX_top,
      SYNC_RST_UART_CLK,
      TX_busy,
      RX_out_valid_top;

wire  I_clk_en_top;

wire  Gate_EN;

wire  [`WIDTH-1:0]  sync_RX_OUT_DATA;
wire  sync_RX_OUT_V;

wire  [`WIDTH-1:0]  CTRL_out_DATA;
wire  CTRL_out_V;

wire  SYNC_TX_busy;
////////////////////////////////////////////////////////////////////////////////
//////////////////////////// internal wires of DFT ////////////////////////////
//////////////////////////////////////////////////////////////////////////////
wire	REF_CLK_M,
	UART_CLK_M,
	CLK_TX_top_M,
	RST_M,
	SYNC_RST_REF_CLK_M,
	SYNC_RST_UART_CLK_M;
////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////// DFT_mux /////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
mux2X1 U0_DFT_MUX_REF_CLK (
	.IN_0(REF_CLK),
	.IN_1(scan_clk),
	.SEL(test_mode),
	.OUT(REF_CLK_M)
);
mux2X1 U0_DFT_MUX_UART_CLK (
	.IN_0(UART_CLK),
	.IN_1(scan_clk),
	.SEL(test_mode),
	.OUT(UART_CLK_M)
);
mux2X1 U0_DFT_MUX_UART_TX_CLK (
	.IN_0(CLK_TX_top),
	.IN_1(scan_clk),
	.SEL(test_mode),
	.OUT(CLK_TX_top_M)
);
mux2X1 U0_DFT_MUX_RST (
	.IN_0(RST),
	.IN_1(scan_rst),
	.SEL(test_mode),
	.OUT(RST_M)
);
mux2X1 U0_DFT_MUX_RST_REF (
	.IN_0(SYNC_RST_REF_CLK),
	.IN_1(scan_rst),
	.SEL(test_mode),
	.OUT(SYNC_RST_REF_CLK_M)
);
mux2X1 U0_DFT_MUX_RST_UART (
	.IN_0(SYNC_RST_UART_CLK),
	.IN_1(scan_rst),
	.SEL(test_mode),
	.OUT(SYNC_RST_UART_CLK_M)
);
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////// SYS_CTRL ////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
SYS_CTRL U0_CTRL_TOP(
    //CTRL_RX
    .UART_RX_DATA(sync_RX_OUT_DATA),
    .UART_RX_VLD(sync_RX_OUT_V),
    .CLK(REF_CLK_M),
    .RST(SYNC_RST_REF_CLK_M),
    .ALU_EN(EN_top),
    .ALU_FUN(ALU_FUN_top),
    .CLKG_EN(Gate_EN),
    .RF_Address(Address_top),
    .RF_WrEn(WrEn_top),
    .RF_RdEn(RdEn_top),
    .RF_WrData(WrData_top),
    //CTRL_TX
    .ALU_OUT(ALU_OUT_top),
    .ALU_OUT_VLD(OUT_VALID_top),
    .RF_RdData(RdData_top),
    .RF_RdData_VLD(RdData_VLD_top),
    .UART_TX_Busy(TX_busy),
    .UART_TX_DATA(CTRL_out_DATA),
    .UART_TX_VLD(CTRL_out_V),
    .CLKDIV_EN(I_clk_en_top)
);
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////// RegFile ////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
RegFile UO_RegFile(
.CLK(REF_CLK_M),
.RST(SYNC_RST_REF_CLK_M),
.WrEn(WrEn_top),
.RdEn(RdEn_top),
.Address(Address_top),
.WrData(WrData_top),
.RdData(RdData_top),
.RdData_VLD(RdData_VLD_top),
.REG0(REG0_OP_A),
.REG1(REG1_OP_B),
.REG2(REG2_UART_convig),
.REG3(REG3_div)
);
////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////// ALU //////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
ALU U0_ALU
(
  .A(REG0_OP_A), 
  .B(REG1_OP_B),
  .EN(EN_top),
  .ALU_FUN(ALU_FUN_top),
  .CLK(ALU_CLK),
  .RST(SYNC_RST_REF_CLK_M),  
  .ALU_OUT(ALU_OUT_top),
  .OUT_VALID(OUT_VALID_top)  
);
////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////// UART /////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
UART_TOP U0_UART(
    .TX_IN_DATA(TX_IN_DATA_top),
    .RX_IN_DATA(RX_IN),
    .TX_IN_valid(TX_IN_valid_top),
    .CLK_RX(UART_CLK_M),
    .CLK_TX(CLK_TX_top_M),
    .parity_enable(REG2_UART_convig[0]),
    .RST(SYNC_RST_UART_CLK_M),
    .parity_type(REG2_UART_convig[1]),
    .prescale(REG2_UART_convig[6:2]),
    .TX_out_valid(TX_busy),
    .RX_out_valid(RX_out_valid_top),
    .TX_out_DATA(TX_OUT),
    .RX_out_DATA(RX_out_DATA_top)
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// clock divider ///////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
clock_divider U0_clock_divider(
  .I_div_ratio(REG3_div[4:0]),     ////////////////////////////////////////
  .I_ref_clk(UART_CLK_M),
  .I_clk_en(I_clk_en_top),
  .I_rst_n(SYNC_RST_UART_CLK_M),
  .o_div_clk(CLK_TX_top) 
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// clock Gating ///////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
CLK_GATE U0_CLK_GATE (
.CLK_EN(Gate_EN || test_mode),
.CLK(REF_CLK_M),
.GATED_CLK(ALU_CLK)
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// Data Sync of RX /////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
data_synchronizer U0_Data_Sync_of_RX (
    .unsync_bus(RX_out_DATA_top),
    .bus_enable(RX_out_valid_top),
    .clk(REF_CLK_M),
    .rst(SYNC_RST_REF_CLK_M),
    .sync_bus(sync_RX_OUT_DATA),
    .enable_pulse(sync_RX_OUT_V)  
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// Data Sync of TX /////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
data_synchronizer U0_Data_Sync_of_TX (
    .unsync_bus(CTRL_out_DATA),
    .bus_enable(CTRL_out_V),
    .clk(CLK_TX_top_M),
    .rst(SYNC_RST_UART_CLK_M),
    .sync_bus(TX_IN_DATA_top),
    .enable_pulse(TX_IN_valid_top)  
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// SYNC RST UART CLK ///////////////////////////////
//////////////////////////////////////////////////////////////////////////////
RST_synchronizer U0_SYNC_RST_UART_CLK (
    .RST(RST_M),
    .clk(UART_CLK_M),
    .SYNC_RST(SYNC_RST_UART_CLK)
);
////////////////////////////////////////////////////////////////////////////////
///////////////////////////// SYNC RST REF CLK ///////////////////////////////
//////////////////////////////////////////////////////////////////////////////
RST_synchronizer U0_SYNC_RST_REF_CLK (
    .RST(RST_M),
    .clk(REF_CLK_M),
    .SYNC_RST(SYNC_RST_REF_CLK)
);
////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////// SYNC Bit //////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
bit_synchronizer U0_bit_synchronizer (
    .ASYNC(TX_busy),
    .RST(SYNC_RST_REF_CLK_M),
    .clk(REF_CLK_M),
    .SYNC(SYNC_TX_busy)
);
endmodule
